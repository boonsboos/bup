module main

import editor

fn main() {
	
	// register plugins here

	// start bup
	editor.start()
}